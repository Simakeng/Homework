EX2                 ;标题
VS 1 0 10           ;电源10V，连接在节点1和节点0
R1 1 2 20           ;电阻R1，20欧姆,连接在节点1和节点2
R2 2 0 20           ;电阻R2，20欧姆,连接在节点2和节点0
R3 3 0 4K           ;电阻R3，4k欧姆,连接在节点3和节点0
L 2 3 0.2 IC=0.2    ;电感L，0.2H,连接在节点2和节点3
C 3 0 0.5U IC=2     ;电容C，0.5微法,连接在节点3和节点0
.TRAN 0.1M 30M UIC  ;瞬态分析,打印时间间隔0.1ms，终止时间30ms，使用初始化条件
.END                ;结束